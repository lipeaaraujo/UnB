CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 212 386 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 TF
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4595 0 0
2
45063 0
0
13 Logic Switch~
5 212 347 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 TD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9395 0 0
2
45063 1
0
7 Ground~
168 621 255 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3303 0 0
2
5.90077e-315 0
0
2 +V
167 217 193 0 1 3
0 3
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4498 0 0
2
5.90077e-315 0
0
7 Ground~
168 617 505 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9728 0 0
2
45063 2
0
9 Inverter~
13 328 450 0 2 22
0 4 8
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3789 0 0
2
45063 3
0
9 Inverter~
13 328 494 0 2 22
0 5 9
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3978 0 0
2
45063 4
0
7 Ground~
168 620 380 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3494 0 0
2
45063 5
0
4 LED~
171 617 484 0 2 2
10 6 2
0
0 0 880 0
4 LED1
17 0 45 8
3 CH3
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3507 0 0
2
45063 6
0
4 LED~
171 620 361 0 2 2
10 7 2
0
0 0 880 0
4 LED1
17 0 45 8
3 CH2
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5151 0 0
2
45063 7
0
4 LED~
171 621 223 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
3 CH1
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3701 0 0
2
45063 8
0
9 Inverter~
13 357 347 0 2 22
0 4 7
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
8585 0 0
2
45063 9
0
9 2-In AND~
219 409 459 0 3 22
0 8 9 6
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8809 0 0
2
45063 10
0
12
2 1 2 0 0 4224 0 11 3 0 0 2
621 233
621 249
1 1 3 0 0 4224 0 4 11 0 0 3
217 202
621 202
621 213
0 1 4 0 0 4096 0 0 6 12 0 3
268 347
268 450
313 450
1 1 5 0 0 4224 0 1 7 0 0 3
224 386
224 494
313 494
3 1 6 0 0 4224 0 13 9 0 0 3
430 459
617 459
617 474
2 1 7 0 0 4224 0 12 10 0 0 3
378 347
620 347
620 351
2 1 8 0 0 4224 0 6 13 0 0 2
349 450
385 450
2 2 9 0 0 8320 0 7 13 0 0 4
349 494
364 494
364 468
385 468
2 1 2 0 0 0 0 10 8 0 0 2
620 371
620 374
1 2 2 0 0 0 0 8 10 0 0 2
620 374
620 371
2 1 2 0 0 0 0 9 5 0 0 2
617 494
617 499
1 1 4 0 0 4224 0 2 12 0 0 2
224 347
342 347
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 201
863 268 1060 452
873 276 1049 420
201 TD TF R  | CH1 CH2 CH3 
0  0  0  | X   X   X 
0  0  1  | X   X   1
0  1  0  | X   1   X
0  1  1  | X   1   0
1  0  0  | 1   X   X
1  0  1  | 1   X   0
1  1  0  | 1   0   X 
1  1  1  | 1   0   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 239
775 106 1172 270
785 114 1161 242
239 Entradas:
A: chave 1 (0: chave fechada, 1: chave aberta)
B: chave 2 (0: chave fechada, 1: chave aberta)
C: chave 3 (0: chave fechada, 1: chave aberta)

Sa�das:
S: detector (0: n�mero de chaves ligadas �mpar,
1: n�mero de chaves par)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 248 102 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45097.7 0
0
13 Logic Switch~
5 226 103 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45097.7 0
0
13 Logic Switch~
5 204 102 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45097.7 0
0
9 3-In AND~
219 446 482 0 4 22
0 15 13 10 2
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
3421 0 0
2
45097.7 0
0
9 3-In AND~
219 446 439 0 4 22
0 14 13 10 3
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
8157 0 0
2
45097.7 0
0
9 3-In AND~
219 446 396 0 4 22
0 15 12 10 4
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
5572 0 0
2
45097.7 0
0
9 3-In AND~
219 446 355 0 4 22
0 14 12 10 5
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 4 0
1 U
8901 0 0
2
45097.7 0
0
9 3-In AND~
219 447 314 0 4 22
0 15 13 11 6
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
7361 0 0
2
45097.7 0
0
9 3-In AND~
219 447 272 0 4 22
0 14 13 11 7
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 3 0
1 U
4747 0 0
2
45097.7 0
0
9 3-In AND~
219 447 230 0 4 22
0 15 12 11 8
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 3 0
1 U
972 0 0
2
45097.7 0
0
9 3-In AND~
219 447 188 0 4 22
0 14 12 11 9
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
3472 0 0
2
45097.7 0
0
9 Inverter~
13 341 146 0 2 22
0 15 14
0
0 0 112 270
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9998 0 0
2
45097.7 0
0
9 Inverter~
13 316 145 0 2 22
0 13 12
0
0 0 112 270
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3536 0 0
2
45097.7 0
0
9 Inverter~
13 292 145 0 2 22
0 10 11
0
0 0 112 270
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4597 0 0
2
45097.7 0
0
35
4 0 2 0 0 4224 0 4 0 0 0 2
467 482
578 482
4 0 3 0 0 4224 0 5 0 0 0 2
467 439
579 439
4 0 4 0 0 4224 0 6 0 0 0 2
467 396
579 396
4 0 5 0 0 4224 0 7 0 0 0 2
467 355
579 355
4 0 6 0 0 4224 0 8 0 0 0 2
468 314
580 314
4 0 7 0 0 4224 0 9 0 0 0 2
468 272
581 272
4 0 8 0 0 4224 0 10 0 0 0 2
468 230
583 230
4 0 9 0 0 4224 0 11 0 0 0 2
468 188
582 188
0 3 10 0 0 8192 0 0 4 10 0 3
204 448
204 491
422 491
0 3 10 0 0 0 0 0 5 11 0 3
204 404
204 448
422 448
0 3 10 0 0 0 0 0 6 12 0 3
204 363
204 405
422 405
0 3 10 0 0 4224 0 0 7 34 0 3
204 127
204 364
422 364
0 3 11 0 0 8320 0 0 8 14 0 3
295 281
295 323
423 323
0 3 11 0 0 0 0 0 9 21 0 3
295 239
295 281
423 281
0 2 12 0 0 8192 0 0 6 16 0 3
319 355
319 396
422 396
0 2 12 0 0 4224 0 0 7 22 0 3
319 230
319 355
422 355
2 0 13 0 0 4096 0 4 0 0 18 3
422 482
226 482
226 439
0 2 13 0 0 0 0 0 5 20 0 3
226 314
226 439
422 439
2 0 13 0 0 4224 0 9 0 0 20 2
423 272
226 272
0 2 13 0 0 0 0 0 8 35 0 3
226 121
226 314
423 314
0 3 11 0 0 0 0 0 10 30 0 3
295 197
295 239
423 239
0 2 12 0 0 0 0 0 10 31 0 3
319 187
319 230
423 230
0 1 14 0 0 4224 0 0 5 24 0 3
344 346
344 430
422 430
0 1 14 0 0 0 0 0 7 25 0 3
344 262
344 346
422 346
0 1 14 0 0 0 0 0 9 32 0 3
344 179
344 263
423 263
0 1 15 0 0 8192 0 0 4 27 0 3
248 387
248 473
422 473
0 1 15 0 0 0 0 0 6 28 0 3
248 305
248 387
422 387
0 1 15 0 0 8320 0 0 8 29 0 3
248 220
248 305
423 305
1 1 15 0 0 0 0 1 10 0 0 3
248 114
248 221
423 221
2 3 11 0 0 0 0 14 11 0 0 3
295 163
295 197
423 197
2 2 12 0 0 0 0 13 11 0 0 3
319 163
319 188
423 188
2 1 14 0 0 0 0 12 11 0 0 3
344 164
344 179
423 179
1 1 15 0 0 0 0 1 12 0 0 3
248 114
344 114
344 128
1 1 10 0 0 0 0 3 14 0 0 3
204 114
204 127
295 127
1 1 13 0 0 0 0 2 13 0 0 4
226 115
226 121
319 121
319 127
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 75 552 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
45063.4 0
0
13 Logic Switch~
5 77 508 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9442 0 0
2
45063.4 0
0
13 Logic Switch~
5 78 469 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9424 0 0
2
45063.4 0
0
13 Logic Switch~
5 79 429 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 MODO
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9968 0 0
2
45063.4 0
0
4 LED~
171 426 330 0 2 2
10 3 2
0
0 0 864 0
4 LED1
17 0 45 8
2 S2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
9281 0 0
2
45063.4 0
0
9 Inverter~
13 243 338 0 2 22
0 7 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
8464 0 0
2
45063.4 0
0
9 3-In AND~
219 251 232 0 4 22
0 8 7 11 9
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
7168 0 0
2
45063.4 0
0
7 Ground~
168 579 388 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3171 0 0
2
45063.4 0
0
4 LED~
171 433 218 0 2 2
10 4 2
0
0 0 864 0
4 LED1
17 0 45 8
2 S1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4139 0 0
2
45063.4 0
0
8 2-In OR~
219 318 203 0 3 22
0 10 9 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6435 0 0
2
45063.4 0
0
9 Inverter~
13 243 302 0 2 22
0 8 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5283 0 0
2
45063.4 0
0
9 2-In AND~
219 327 320 0 3 22
0 6 5 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6874 0 0
2
45063.4 0
0
9 3-In AND~
219 251 179 0 4 22
0 8 7 12 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
5305 0 0
2
45063.4 0
0
16
2 0 2 0 0 4096 0 5 0 0 3 2
426 340
579 340
3 1 3 0 0 4224 0 12 5 0 0 2
348 320
426 320
2 1 2 0 0 8320 0 9 8 0 0 3
433 228
579 228
579 382
3 1 4 0 0 4224 0 10 9 0 0 3
351 203
433 203
433 208
2 2 5 0 0 12416 0 6 12 0 0 4
264 338
279 338
279 329
303 329
2 1 6 0 0 12416 0 11 12 0 0 4
264 302
279 302
279 311
303 311
1 0 7 0 0 4096 0 6 0 0 14 2
228 338
129 338
1 0 8 0 0 4096 0 11 0 0 16 2
228 302
114 302
4 2 9 0 0 8320 0 7 10 0 0 4
272 232
291 232
291 212
305 212
4 1 10 0 0 4224 0 13 10 0 0 4
272 179
291 179
291 194
305 194
1 3 11 0 0 8320 0 1 7 0 0 4
87 552
161 552
161 241
227 241
1 3 12 0 0 8320 0 2 13 0 0 4
89 508
145 508
145 188
227 188
2 0 7 0 0 0 0 7 0 0 14 2
227 232
129 232
1 2 7 0 0 8320 0 3 13 0 0 4
90 469
129 469
129 179
227 179
1 0 8 0 0 0 0 7 0 0 16 2
227 223
114 223
1 1 8 0 0 8320 0 4 13 0 0 4
91 429
114 429
114 170
227 170
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 373
848 211 1037 555
858 219 1026 491
373 MODO A  B  C  | S1 S2
0    0  0  0  | 0  1
0    0  0  1  | 0  1
0    0  1  0  | 0  1
0    0  1  1  | 0  1
0    1  0  0  | 0  0
0    1  0  1  | 0  0
0    1  1  0  | 0  0
0    1  1  1  | 0  0
1    0  0  0  | 0  0
1    0  0  1  | 0  0
1    0  1  0  | 0  0
1    0  1  1  | 0  0
1    1  0  0  | 0  0
1    1  0  1  | 1  0
1    1  1  0  | 1  0
1    1  1  1  | 1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 337
617 28 1166 212
627 36 1155 180
337 Entradas:
MODO: bot�o MODO (0: bot�o n�o acionado, 1: bot�o acionado)
A, B e C: indicam o valor de combust�vel presente no tanque de 
combust�vel, com 000 representado tanque vazio e 111 representando 
tanque cheio.

Sa�das:
S1: sinal da luz verde, (0: desligada, 1: ligada)
S2: sinal da luz vermelha, (0: desligada, 1: ligada)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

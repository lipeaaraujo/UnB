CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 511 166 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 492 166 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 452 166 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 435 166 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 399 166 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 378 166 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 338 166 0 1 11
0 33
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.90081e-315 0
0
13 Logic Switch~
5 316 166 0 1 11
0 34
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90081e-315 0
0
9 4-In AND~
219 457 597 0 5 22
0 6 7 8 9 3
0
0 0 112 270
6 74LS21
-21 -28 21 -20
3 U9A
19 -4 40 4
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 9 0
1 U
4747 0 0
2
5.90081e-315 0
0
8 4-In OR~
219 601 592 0 5 22
0 13 12 11 10 4
0
0 0 112 270
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
972 0 0
2
5.90081e-315 0
0
8 4-In OR~
219 305 594 0 5 22
0 17 18 19 20 5
0
0 0 112 270
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3472 0 0
2
5.90081e-315 0
0
7 Ground~
168 803 702 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
5.90081e-315 0
0
4 LED~
171 604 653 0 2 2
10 4 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3536 0 0
2
5.90081e-315 0
0
4 LED~
171 455 651 0 2 2
10 3 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4597 0 0
2
5.90081e-315 0
0
4 LED~
171 308 653 0 2 2
10 5 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3835 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 619 488 0 3 22
0 14 7 13
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U7B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3670 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 514 489 0 3 22
0 15 8 12
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U7A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5616 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 410 486 0 3 22
0 16 9 11
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U5D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 570 489 0 3 22
0 21 7 17
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
317 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 464 488 0 3 22
0 22 8 18
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3108 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 363 486 0 3 22
0 23 9 19
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 598 390 0 3 22
0 26 25 21
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
5.90081e-315 5.30499e-315
0
9 Inverter~
13 626 391 0 2 22
0 26 6
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U3D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
7876 0 0
2
5.90081e-315 5.26354e-315
0
9 2-In AND~
219 661 390 0 3 22
0 24 26 14
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6369 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 499 384 0 3 22
0 27 29 22
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9172 0 0
2
5.90081e-315 5.30499e-315
0
9 Inverter~
13 527 385 0 2 22
0 27 7
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U3C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
7100 0 0
2
5.90081e-315 5.26354e-315
0
9 2-In AND~
219 562 384 0 3 22
0 28 27 15
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3820 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 394 390 0 3 22
0 32 31 23
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7678 0 0
2
5.90081e-315 5.30499e-315
0
9 Inverter~
13 422 391 0 2 22
0 32 8
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U3B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
961 0 0
2
5.90081e-315 5.26354e-315
0
9 2-In AND~
219 457 390 0 3 22
0 30 32 16
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3178 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 359 390 0 3 22
0 33 35 10
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3409 0 0
2
5.90081e-315 0
0
9 Inverter~
13 324 391 0 2 22
0 35 9
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3951 0 0
2
5.90081e-315 0
0
9 2-In AND~
219 296 390 0 3 22
0 35 34 20
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8885 0 0
2
5.90081e-315 0
0
9 2-In XOR~
219 626 295 0 3 22
0 24 25 26
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U1D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3780 0 0
2
5.90081e-315 0
0
9 2-In XOR~
219 527 294 0 3 22
0 28 29 27
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U1C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9265 0 0
2
5.90081e-315 0
0
9 2-In XOR~
219 422 296 0 3 22
0 30 31 32
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U1B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9442 0 0
2
5.90081e-315 0
0
9 2-In XOR~
219 324 295 0 3 22
0 33 34 35
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U1A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9424 0 0
2
5.90081e-315 0
0
61
5 1 3 0 0 4224 0 9 14 0 0 2
455 620
455 641
5 0 4 0 0 0 0 10 0 0 7 2
604 622
604 622
5 0 5 0 0 0 0 11 0 0 8 2
308 624
308 624
2 0 2 0 0 8192 0 15 0 0 5 3
308 663
308 687
455 687
2 0 2 0 0 8192 0 14 0 0 6 3
455 661
455 687
604 687
2 1 2 0 0 8320 0 13 12 0 0 4
604 663
604 687
803 687
803 696
0 1 4 0 0 4224 0 0 13 0 0 2
604 618
604 643
0 1 5 0 0 4224 0 0 15 0 0 2
308 620
308 643
2 1 6 0 0 16512 0 23 9 0 0 6
629 409
629 456
637 456
637 557
468 557
468 575
0 2 7 0 0 4224 0 0 9 28 0 4
530 458
530 553
459 553
459 575
0 3 8 0 0 4224 0 0 9 30 0 4
425 458
425 553
450 553
450 575
0 4 9 0 0 8320 0 0 9 32 0 4
327 457
327 557
441 557
441 575
3 4 10 0 0 12416 0 31 10 0 0 5
357 413
381 413
381 541
590 541
590 572
3 3 11 0 0 8320 0 18 10 0 0 4
408 509
408 530
599 530
599 572
3 2 12 0 0 8320 0 17 10 0 0 4
512 512
512 520
608 520
608 572
3 1 13 0 0 4224 0 16 10 0 0 2
617 511
617 572
3 1 14 0 0 8320 0 24 16 0 0 4
659 413
659 438
626 438
626 466
0 2 7 0 0 0 0 0 16 28 0 3
530 449
608 449
608 466
3 1 15 0 0 8320 0 27 17 0 0 4
560 407
560 439
521 439
521 467
0 2 8 0 0 0 0 0 17 30 0 3
425 449
503 449
503 467
3 1 16 0 0 8320 0 30 18 0 0 4
455 413
455 439
417 439
417 464
0 2 9 0 0 0 0 0 18 32 0 3
327 439
399 439
399 464
3 1 17 0 0 8320 0 19 11 0 0 4
568 512
568 546
321 546
321 574
3 2 18 0 0 8320 0 20 11 0 0 4
462 511
462 536
312 536
312 574
3 3 19 0 0 8320 0 21 11 0 0 4
361 509
361 528
303 528
303 574
3 4 20 0 0 4224 0 33 11 0 0 2
294 413
294 574
3 1 21 0 0 4224 0 22 19 0 0 4
596 413
596 458
577 458
577 467
2 2 7 0 0 0 0 26 19 0 0 4
530 403
530 458
559 458
559 467
3 1 22 0 0 4224 0 25 20 0 0 4
497 407
497 458
471 458
471 466
2 2 8 0 0 0 0 29 20 0 0 4
425 409
425 458
453 458
453 466
3 1 23 0 0 4224 0 28 21 0 0 4
392 413
392 458
370 458
370 464
2 2 9 0 0 0 0 32 21 0 0 4
327 409
327 458
352 458
352 464
0 1 24 0 0 8192 0 0 24 54 0 3
638 272
668 272
668 368
0 2 25 0 0 8192 0 0 22 55 0 3
620 272
587 272
587 368
0 1 26 0 0 4096 0 0 22 36 0 3
629 358
605 358
605 368
0 2 26 0 0 0 0 0 24 37 0 3
629 358
650 358
650 368
3 1 26 0 0 4224 0 34 23 0 0 2
629 325
629 373
3 0 27 0 0 0 0 35 0 0 43 2
530 324
530 324
0 1 28 0 0 8320 0 0 27 56 0 3
539 266
569 266
569 362
0 2 29 0 0 8320 0 0 25 57 0 3
521 266
488 266
488 362
0 1 27 0 0 4096 0 0 25 42 0 3
530 352
506 352
506 362
0 2 27 0 0 0 0 0 27 43 0 3
530 352
551 352
551 362
3 1 27 0 0 4224 0 0 26 0 0 2
530 319
530 367
0 1 30 0 0 8320 0 0 30 60 0 3
434 272
464 272
464 368
0 2 31 0 0 8320 0 0 28 61 0 3
416 272
383 272
383 368
0 1 32 0 0 4096 0 0 28 47 0 3
425 358
401 358
401 368
0 2 32 0 0 0 0 0 30 48 0 3
425 358
446 358
446 368
3 1 32 0 0 4224 0 36 29 0 0 2
425 326
425 373
0 1 33 0 0 8320 0 0 31 58 0 3
338 272
366 272
366 368
0 2 34 0 0 8320 0 0 33 59 0 3
316 272
285 272
285 368
0 1 35 0 0 4096 0 0 33 52 0 3
327 358
303 358
303 368
0 2 35 0 0 0 0 0 31 53 0 3
327 358
348 358
348 368
3 1 35 0 0 4224 0 37 32 0 0 2
327 325
327 373
1 1 24 0 0 8320 0 1 34 0 0 4
511 178
511 195
638 195
638 276
1 2 25 0 0 8320 0 2 34 0 0 4
492 178
492 203
620 203
620 276
1 1 28 0 0 0 0 3 35 0 0 4
452 178
452 226
539 226
539 275
1 2 29 0 0 0 0 4 35 0 0 4
435 178
435 236
521 236
521 275
1 1 33 0 0 0 0 7 37 0 0 4
338 178
338 272
336 272
336 276
1 2 34 0 0 0 0 8 37 0 0 4
316 178
316 272
318 272
318 276
1 1 30 0 0 0 0 5 36 0 0 4
399 178
399 255
434 255
434 277
1 2 31 0 0 0 0 6 36 0 0 4
378 178
378 263
416 263
416 277
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 71 269 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 S
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 72 226 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90077e-315 0
0
9 Inverter~
13 190 334 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3124 0 0
2
5.90077e-315 0
0
4 LED~
171 440 359 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 E2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3421 0 0
2
5.90077e-315 0
0
7 Ground~
168 440 418 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
5.90077e-315 0
0
9 Inverter~
13 190 274 0 2 22
0 5 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
5572 0 0
2
5.90077e-315 0
0
9 2-In AND~
219 296 265 0 3 22
0 4 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
5.90077e-315 0
0
4 LED~
171 440 304 0 2 2
10 6 3
0
0 0 880 0
4 LED1
17 0 45 8
2 E1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
5.90077e-315 0
0
8
2 0 3 0 0 8320 0 3 0 0 3 2
211 334
440 334
0 1 4 0 0 4096 0 0 3 5 0 3
137 226
137 334
175 334
2 1 3 0 0 16 0 8 4 0 0 2
440 314
440 349
2 1 2 0 0 4224 0 4 5 0 0 2
440 369
440 412
1 1 4 0 0 4224 0 2 7 0 0 4
84 226
255 226
255 256
272 256
1 1 5 0 0 4224 0 1 6 0 0 4
83 269
157 269
157 274
175 274
3 1 6 0 0 4224 0 7 8 0 0 3
317 265
440 265
440 294
2 2 7 0 0 4224 0 6 7 0 0 2
211 274
272 274
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 69
743 317 868 421
753 325 857 405
69 B S | E1 | E2
0 0 | 0  | 1
0 1 | 0  | 1
1 0 | 1  | 0
1 1 | 0  | 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 266
614 136 1059 300
624 144 1048 272
266 Entradas:
B: bot�o, (0: bot�o desligado, 1: bot�o ligado)
S: sensor de n�vel m�ximo, (0: n�vel m�ximo n�o 
atingido, 1: n�vel m�ximo atingido).

Sa�das:
E1: Eletrov�lvula de entrada, (0: fechada, 1: aberta)
E2: Eletrov�lvula de sa�da, (0: fechada, 1: aberta)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

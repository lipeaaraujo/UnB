CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 111 258 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45114.8 0
0
13 Logic Switch~
5 112 214 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45114.8 0
0
8 2-In OR~
219 639 360 0 3 22
0 7 6 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3124 0 0
2
45114.8 0
0
9 2-In AND~
219 599 337 0 3 22
0 5 4 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3421 0 0
2
45114.8 0
0
9 2-In AND~
219 599 383 0 3 22
0 3 2 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8157 0 0
2
45114.8 0
0
8 3-In OR~
219 647 488 0 4 22
0 9 10 11 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
5572 0 0
2
45114.8 0
0
5 7415~
219 599 443 0 4 22
0 12 5 4 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 4 0
1 U
8901 0 0
2
45114.8 0
0
5 7415~
219 599 489 0 4 22
0 4 2 13 10
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
7361 0 0
2
45114.8 0
0
5 7415~
219 598 533 0 4 22
0 3 2 12 11
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
4747 0 0
2
45114.8 0
0
8 2-In OR~
219 613 620 0 3 22
0 13 5 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
972 0 0
2
45114.8 0
0
9 2-In AND~
219 610 740 0 3 22
0 13 2 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3472 0 0
2
45114.8 0
0
2 +V
167 571 276 0 1 3
0 17
0
0 0 54256 90
2 5V
-8 -15 6 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
45114.8 0
0
9 Inverter~
13 206 314 0 2 22
0 20 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3536 0 0
2
45114.8 0
0
6 74LS73
102 316 323 0 12 25
0 14 15 19 18 8 17 19 18 3
4 13 12
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 0 0 0 0 0
1 U
4597 0 0
2
45114.8 0
0
7 74LS175
131 315 216 0 14 29
0 18 20 21 22 23 16 24 25 26
27 28 29 2 5
0
0 0 4848 0
6 74F175
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3835 0 0
2
45114.8 0
0
44
0 2 2 0 0 8192 0 0 5 37 0 3
533 394
533 392
575 392
0 1 3 0 0 8192 0 0 5 35 0 3
517 373
517 374
575 374
0 2 4 0 0 4096 0 0 4 34 0 2
509 346
575 346
0 1 5 0 0 8192 0 0 4 36 0 3
525 327
525 328
575 328
3 2 6 0 0 4224 0 5 3 0 0 3
620 383
620 369
626 369
3 1 7 0 0 4224 0 4 3 0 0 3
620 337
620 351
626 351
3 0 8 0 0 4096 0 3 0 0 30 2
672 360
686 360
4 1 9 0 0 4224 0 7 6 0 0 3
620 443
620 479
634 479
4 2 10 0 0 8320 0 8 6 0 0 3
620 489
620 488
635 488
4 3 11 0 0 4224 0 9 6 0 0 3
619 533
619 497
634 497
0 1 3 0 0 0 0 0 9 35 0 3
517 523
517 524
574 524
0 2 2 0 0 0 0 0 9 37 0 3
533 532
533 533
574 533
0 3 12 0 0 4096 0 0 9 32 0 2
542 542
574 542
0 3 13 0 0 4096 0 0 8 33 0 2
552 498
575 498
0 2 2 0 0 0 0 0 8 37 0 3
533 488
533 489
575 489
0 1 4 0 0 0 0 0 8 34 0 3
509 478
509 480
575 480
0 3 4 0 0 0 0 0 7 34 0 3
509 451
509 452
575 452
0 2 5 0 0 0 0 0 7 36 0 2
525 443
575 443
0 1 12 0 0 4096 0 0 7 32 0 2
542 434
575 434
0 2 5 0 0 8192 0 0 10 36 0 3
525 628
525 629
600 629
0 1 13 0 0 8192 0 0 10 33 0 3
552 610
552 611
600 611
0 0 3 0 0 8192 0 0 0 35 0 3
517 821
407 821
407 509
0 0 2 0 0 8192 0 0 0 37 0 3
533 810
419 810
419 510
0 0 13 0 0 8192 0 0 0 33 0 3
552 801
430 801
430 508
3 1 14 0 0 8320 0 11 14 0 0 8
631 740
724 740
724 115
203 115
203 279
265 279
265 296
284 296
0 2 2 0 0 0 0 0 11 37 0 3
533 747
533 749
586 749
0 1 13 0 0 0 0 0 11 33 0 3
552 728
552 731
586 731
3 2 15 0 0 16512 0 10 14 0 0 9
646 620
646 622
712 622
712 128
212 128
212 289
253 289
253 305
284 305
4 6 16 0 0 16512 0 6 15 0 0 7
680 488
680 507
698 507
698 140
219 140
219 243
283 243
0 5 8 0 0 8336 0 0 14 0 0 5
686 421
686 150
226 150
226 332
284 332
1 6 17 0 0 8320 0 12 14 0 0 5
582 274
582 158
235 158
235 341
284 341
12 0 12 0 0 8320 0 14 0 0 0 3
354 350
542 350
542 849
11 0 13 0 0 8320 0 14 0 0 0 3
348 341
552 341
552 859
10 0 4 0 0 8320 0 14 0 0 0 3
354 314
509 314
509 858
9 0 3 0 0 8320 0 14 0 0 0 3
348 305
517 305
517 862
14 0 5 0 0 8320 0 15 0 0 0 3
353 252
525 252
525 856
13 0 2 0 0 8320 0 15 0 0 0 3
347 243
533 243
533 847
0 8 18 0 0 8192 0 0 14 39 0 3
245 328
245 359
278 359
0 4 18 0 0 4096 0 0 14 43 0 5
179 258
179 328
245 328
245 323
278 323
0 7 19 0 0 4096 0 0 14 41 0 3
261 314
261 350
278 350
2 3 19 0 0 4224 0 13 14 0 0 2
227 314
278 314
0 1 20 0 0 4096 0 0 13 44 0 3
140 212
140 314
191 314
1 1 18 0 0 12416 0 1 15 0 0 4
123 258
180 258
180 189
277 189
2 1 20 0 0 4224 0 15 2 0 0 4
283 198
140 198
140 214
124 214
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

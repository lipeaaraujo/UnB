CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 79 829 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 P
-3 -25 4 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
45063.8 0
0
13 Logic Switch~
5 78 901 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3409 0 0
2
45063.8 7
0
13 Logic Switch~
5 77 939 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
45063.8 2
0
13 Logic Switch~
5 77 978 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 C1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
45063.8 1
0
13 Logic Switch~
5 77 1015 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
45063.8 0
0
13 Logic Switch~
5 116 365 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9265 0 0
2
45063.8 0
0
13 Logic Switch~
5 116 328 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9442 0 0
2
45063.8 0
0
13 Logic Switch~
5 116 289 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9424 0 0
2
45063.8 0
0
13 Logic Switch~
5 117 251 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -25 4 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9968 0 0
2
45063.8 0
0
6 74266~
219 417 891 0 3 22
0 5 4 3
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9281 0 0
2
45063.8 0
0
4 LED~
171 582 930 0 2 2
10 3 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8464 0 0
2
45063.8 0
0
6 74136~
219 177 920 0 3 22
0 11 10 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7168 0 0
2
45063.8 6
0
6 74136~
219 177 995 0 3 22
0 9 8 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3171 0 0
2
45063.8 5
0
6 74136~
219 262 954 0 3 22
0 6 7 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4139 0 0
2
45063.8 4
0
7 Ground~
168 582 977 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6435 0 0
2
45063.8 3
0
7 Ground~
168 453 353 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5283 0 0
2
45063.8 0
0
6 74136~
219 301 304 0 3 22
0 13 14 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6874 0 0
2
45063.8 0
0
6 74136~
219 216 345 0 3 22
0 16 15 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5305 0 0
2
45063.8 0
0
6 74136~
219 216 270 0 3 22
0 18 17 13
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
34 0 0
2
45063.8 0
0
4 LED~
171 453 319 0 2 2
10 12 2
0
0 0 864 0
4 LED1
17 0 45 8
1 P
27 -10 34 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
969 0 0
2
45063.8 0
0
18
3 1 3 0 0 4224 0 10 11 0 0 3
456 891
582 891
582 920
3 2 4 0 0 4224 0 14 10 0 0 4
295 954
352 954
352 900
401 900
1 1 5 0 0 4224 0 1 10 0 0 4
91 829
352 829
352 882
401 882
2 1 2 0 0 4224 0 11 15 0 0 2
582 940
582 971
3 1 6 0 0 8320 0 12 14 0 0 3
210 920
210 945
246 945
3 2 7 0 0 8320 0 13 14 0 0 3
210 995
210 963
246 963
1 2 8 0 0 4224 0 5 13 0 0 4
89 1015
149 1015
149 1004
161 1004
1 1 9 0 0 4224 0 4 13 0 0 4
89 978
149 978
149 986
161 986
1 2 10 0 0 4224 0 3 12 0 0 4
89 939
149 939
149 929
161 929
1 1 11 0 0 4224 0 2 12 0 0 4
90 901
149 901
149 911
161 911
2 1 2 0 0 0 0 20 16 0 0 2
453 329
453 347
3 1 12 0 0 4224 0 17 20 0 0 3
334 304
453 304
453 309
3 1 13 0 0 8320 0 19 17 0 0 3
249 270
249 295
285 295
3 2 14 0 0 8320 0 18 17 0 0 3
249 345
249 313
285 313
1 2 15 0 0 4224 0 6 18 0 0 4
128 365
188 365
188 354
200 354
1 1 16 0 0 4224 0 7 18 0 0 4
128 328
188 328
188 336
200 336
1 2 17 0 0 4224 0 8 19 0 0 4
128 289
188 289
188 279
200 279
1 1 18 0 0 4224 0 9 19 0 0 4
129 251
188 251
188 261
200 261
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
303 954 340 978
313 962 329 978
2 P1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 65
793 817 894 941
803 825 883 921
65 P  P1  | V
0  0   | 1
0  1   | 0      
1  0   | 0
1  1   | 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 366
550 614 1115 818
560 622 1104 782
366 Entradas:
P: bit de paridade recebido, (0: n�mero par de bits de valor "1", 1: 
n�mero �mpar de bits de valor "1")
A1, B1, C1 e D1: bits de informa��o do transmissor recebidos, s�o 
usados para calcular um segundo bit de paridade P1, que � comparado 
com P.

Sa�das:
V: sinal de verifica��o, (0: bits de paridade diferentes, 1: bits de 
paridade iguais)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 287
726 130 867 474
736 138 856 410
287 A  B  C  D  | P
0  0  0  0  | 0
0  0  0  1  | 1
0  0  1  0  | 1
0  0  1  1  | 0
0  1  0  0  | 1
0  1  0  1  | 0
0  1  1  0  | 0
0  1  1  1  | 1
1  0  0  0  | 1
1  0  0  1  | 0
1  0  1  0  | 0
1  0  1  1  | 1
1  1  0  0  | 0
1  1  0  1  | 1
1  1  1  0  | 1
1  1  1  1  | 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 196
516 13 1089 137
526 21 1078 117
196 Entradas:
A, B, C e D: representam os bits da informa��o do transmissor.

Sa�das:
P: representa o bit de paridade, (0: n�mero par de bits de valor "1", 
1: n�mero �mpar de bits de valor "1")
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
470 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 124 620 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 125 579 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3674 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 125 538 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5697 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 125 496 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3805 0 0
2
5.90077e-315 0
0
9 3-In AND~
219 341 557 0 4 22
0 6 7 8 4
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 8 0
1 U
5219 0 0
2
5.90077e-315 0
0
9 Inverter~
13 245 590 0 2 22
0 9 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3795 0 0
2
5.90077e-315 0
0
9 Inverter~
13 246 557 0 2 22
0 10 7
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3637 0 0
2
5.90077e-315 0
0
9 Inverter~
13 247 523 0 2 22
0 11 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3226 0 0
2
5.90077e-315 0
0
9 Inverter~
13 248 492 0 2 22
0 12 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
6966 0 0
2
5.90077e-315 0
0
9 Inverter~
13 253 421 0 2 22
0 11 17
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9796 0 0
2
5.90077e-315 0
0
9 Inverter~
13 254 333 0 2 22
0 10 18
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
5952 0 0
2
5.90077e-315 0
0
9 3-In AND~
219 322 421 0 4 22
0 12 17 10 16
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 5 0
1 U
3649 0 0
2
5.90077e-315 0
0
9 3-In AND~
219 323 333 0 4 22
0 12 18 9 15
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
3716 0 0
2
5.90077e-315 0
0
8 3-In OR~
219 434 333 0 4 22
0 14 15 16 13
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
4797 0 0
2
5.90077e-315 0
0
9 3-In AND~
219 323 257 0 4 22
0 12 11 19 14
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
4681 0 0
2
5.90077e-315 0
0
9 4-In AND~
219 312 105 0 5 22
0 12 11 10 9 20
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
9730 0 0
2
5.90077e-315 0
0
4 LED~
171 556 527 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 S3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9874 0 0
2
5.90077e-315 0
0
4 LED~
171 556 343 0 2 2
10 13 2
0
0 0 880 0
4 LED1
17 0 45 8
2 S2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
364 0 0
2
5.90077e-315 0
0
9 Inverter~
13 253 281 0 2 22
0 9 19
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3656 0 0
2
5.90077e-315 0
0
8 2-In OR~
219 413 517 0 3 22
0 5 4 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3131 0 0
2
5.90077e-315 0
0
4 LED~
171 561 134 0 2 2
10 20 2
0
0 0 880 0
4 LED1
17 0 45 8
2 S1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6772 0 0
2
5.90077e-315 0
0
7 Ground~
168 843 615 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9557 0 0
2
5.90077e-315 0
0
34
2 0 2 0 0 4096 0 17 0 0 34 2
556 537
843 537
3 1 3 0 0 4224 0 20 17 0 0 2
446 517
556 517
4 2 4 0 0 8320 0 5 20 0 0 4
362 557
378 557
378 526
400 526
2 1 5 0 0 4224 0 9 20 0 0 4
269 492
378 492
378 508
400 508
2 1 6 0 0 4224 0 8 5 0 0 4
268 523
294 523
294 548
317 548
2 2 7 0 0 4224 0 7 5 0 0 2
267 557
317 557
2 3 8 0 0 4224 0 6 5 0 0 4
266 590
294 590
294 566
317 566
1 0 9 0 0 4096 0 6 0 0 30 2
230 590
186 590
1 0 10 0 0 4096 0 7 0 0 31 2
231 557
173 557
1 0 11 0 0 4096 0 8 0 0 32 2
232 523
163 523
1 0 12 0 0 4096 0 9 0 0 33 2
233 492
153 492
2 0 2 0 0 0 0 18 0 0 34 2
556 353
843 353
4 1 13 0 0 4224 0 14 18 0 0 2
467 333
556 333
4 1 14 0 0 8320 0 15 14 0 0 4
344 257
376 257
376 324
421 324
4 2 15 0 0 4224 0 13 14 0 0 2
344 333
422 333
4 3 16 0 0 8320 0 12 14 0 0 4
343 421
376 421
376 342
421 342
0 3 10 0 0 4096 0 0 12 31 0 4
173 444
282 444
282 430
298 430
2 2 17 0 0 4224 0 10 12 0 0 2
274 421
298 421
0 1 11 0 0 4096 0 0 10 32 0 2
163 421
238 421
0 3 9 0 0 4096 0 0 13 30 0 4
186 353
281 353
281 342
299 342
2 2 18 0 0 4224 0 11 13 0 0 2
275 333
299 333
0 1 10 0 0 0 0 0 11 31 0 2
173 333
239 333
2 0 11 0 0 4096 0 15 0 0 32 2
299 257
163 257
2 3 19 0 0 12416 0 19 15 0 0 4
274 281
281 281
281 266
299 266
0 1 9 0 0 0 0 0 19 30 0 3
186 277
186 281
238 281
0 1 12 0 0 4096 0 0 12 33 0 4
153 390
281 390
281 412
298 412
0 1 12 0 0 0 0 0 13 33 0 4
153 301
281 301
281 324
299 324
0 1 12 0 0 0 0 0 15 33 0 4
153 234
281 234
281 248
299 248
5 1 20 0 0 4224 0 16 21 0 0 3
333 105
561 105
561 124
1 4 9 0 0 8320 0 1 16 0 0 4
136 620
186 620
186 119
288 119
1 3 10 0 0 8320 0 2 16 0 0 4
137 579
173 579
173 110
288 110
1 2 11 0 0 8320 0 3 16 0 0 4
137 538
163 538
163 101
288 101
1 1 12 0 0 8320 0 4 16 0 0 4
137 496
153 496
153 92
288 92
2 1 2 0 0 8320 0 21 22 0 0 3
561 144
843 144
843 609
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 390
1024 285 1221 629
1034 293 1210 565
390 A  B  C  D  | S1 S2 S3
0  0  0  0  | 0  0  1
0  0  0  1  | 0  0  1
0  0  1  0  | 0  0  1
0  0  1  1  | 0  0  1
0  1  0  0  | 0  0  1
0  1  0  1  | 0  0  1
0  1  1  0  | 0  0  1
0  1  1  1  | 0  0  1
1  0  0  0  | 0  0  1
1  0  0  1  | 0  1  0
1  0  1  0  | 0  1  0
1  0  1  1  | 0  1  0
1  1  0  0  | 0  1  0
1  1  0  1  | 0  1  0
1  1  1  0  | 0  1  0
1  1  1  1  | 1  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 525
912 41 1469 305
922 49 1458 257
525 Entradas:
A: voto do juiz A (0: voto de qualidade contra,
1: voto de qualidade a favor)
B: voto do juiz B (0: voto contra, 1: voto a favor)
C: voto do juiz C (0: voto contra, 1: voto a favor)
D: voto do juiz D (0: voto contra, 1: voto a favor)

Sa�das:
S1: decis�o a favor por unanimidade,
(0: decis�o n�o un�nime ou n�o a favor, 1: decis�o a favor un�nime)
S2: decis�o a favor por maioria,
(0: decis�o un�nime ou contra, 1: decis�o a favor por maioria)
S3: decis�o contra, (0: decis�o a favor, 1: decis�o contra)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

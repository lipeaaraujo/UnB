CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
250 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 280 160 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
45062.9 0
0
13 Logic Switch~
5 279 125 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7804 0 0
2
45062.9 1
0
13 Logic Switch~
5 280 91 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5523 0 0
2
45062.9 2
0
8 3-In OR~
219 595 225 0 4 22
0 4 5 6 3
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
3330 0 0
2
45062.9 3
0
9 Inverter~
13 383 211 0 2 22
0 10 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3465 0 0
2
45062.9 4
0
9 Inverter~
13 383 304 0 2 22
0 8 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8396 0 0
2
45062.9 5
0
9 Inverter~
13 382 418 0 2 22
0 7 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3685 0 0
2
45062.9 6
0
9 3-In AND~
219 469 202 0 4 22
0 8 7 9 4
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 1 0
1 U
7849 0 0
2
45062.9 7
0
9 3-In AND~
219 467 313 0 4 22
0 11 7 10 5
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
6343 0 0
2
45062.9 8
0
9 3-In AND~
219 467 418 0 4 22
0 8 12 10 6
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
7376 0 0
2
45062.9 9
0
7 Ground~
168 898 366 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9156 0 0
2
45062.9 10
0
4 LED~
171 726 242 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5776 0 0
2
45062.9 11
0
17
4 1 3 0 0 4224 0 4 12 0 0 3
628 225
726 225
726 232
4 1 4 0 0 4224 0 8 4 0 0 4
490 202
554 202
554 216
582 216
4 2 5 0 0 8320 0 9 4 0 0 4
488 313
554 313
554 225
583 225
4 3 6 0 0 8320 0 10 4 0 0 4
488 418
565 418
565 234
582 234
0 2 7 0 0 4096 0 0 8 15 0 4
326 184
411 184
411 202
445 202
0 1 8 0 0 4096 0 0 8 16 0 4
338 167
425 167
425 193
445 193
2 3 9 0 0 4224 0 5 8 0 0 2
404 211
445 211
0 1 10 0 0 8192 0 0 5 13 0 3
312 209
312 211
368 211
0 3 10 0 0 4096 0 0 9 13 0 4
312 337
421 337
421 322
443 322
0 2 7 0 0 0 0 0 9 15 0 4
326 323
408 323
408 313
443 313
2 1 11 0 0 4224 0 6 9 0 0 2
404 304
443 304
0 1 8 0 0 0 0 0 6 16 0 2
338 304
368 304
1 3 10 0 0 8320 0 1 10 0 0 6
292 160
312 160
312 438
408 438
408 427
443 427
2 2 12 0 0 4224 0 7 10 0 0 2
403 418
443 418
1 1 7 0 0 8320 0 2 7 0 0 4
291 125
326 125
326 418
367 418
1 1 8 0 0 8320 0 3 10 0 0 6
292 91
338 91
338 393
416 393
416 409
443 409
2 1 2 0 0 8320 0 12 11 0 0 4
726 252
726 254
898 254
898 360
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 124
1049 278 1166 462
1059 286 1155 430
124 A  B  C  | S
0  0  0  | 0
0  0  1  | 0
0  1  0  | 0
0  1  1  | 1
1  0  0  | 0
1  0  1  | 1
1  1  0  | 1
1  1  1  | 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 239
937 119 1334 283
947 127 1323 255
239 Entradas:
A: chave 1 (0: chave fechada, 1: chave aberta)
B: chave 2 (0: chave fechada, 1: chave aberta)
C: chave 3 (0: chave fechada, 1: chave aberta)

Sa�das:
S: detector (0: n�mero de chaves ligadas �mpar,
1: n�mero de chaves par)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 171 298 0 1 11
0 8
0
0 0 21360 0
2 0V
-50 -3 -36 5
3 Cin
-34 -3 -13 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
45097.7 0
0
13 Logic Switch~
5 171 313 0 1 11
0 7
0
0 0 21360 0
2 0V
-44 -3 -30 5
1 A
-22 -3 -15 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
45097.7 0
0
13 Logic Switch~
5 171 328 0 1 11
0 6
0
0 0 21360 0
2 0V
-43 -4 -29 4
1 B
-22 -4 -15 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
45097.7 0
0
7 Ground~
168 655 370 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9323 0 0
2
45097.7 0
0
4 LED~
171 642 320 0 2 2
10 3 2
0
0 0 352 90
4 Cout
20 -2 48 6
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
317 0 0
2
45097.7 0
0
4 LED~
171 642 294 0 2 2
10 5 2
0
0 0 352 90
1 S
17 -2 24 6
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3108 0 0
2
45097.7 0
0
7 74LS151
20 289 428 0 14 29
0 4 4 4 2 4 2 2 2 2
8 7 6 3 9
0
0 0 4848 512
7 74LS151
-24 -60 25 -52
2 U2
-2 -61 12 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
4299 0 0
2
45097.7 0
0
7 Ground~
168 400 100 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9672 0 0
2
45097.7 0
0
7 Ground~
168 234 103 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7876 0 0
2
45097.7 0
0
2 +V
167 368 101 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6369 0 0
2
45097.7 0
0
7 74LS151
20 291 220 0 14 29
0 4 2 2 4 2 4 4 2 2
8 7 6 5 10
0
0 0 4848 512
7 74LS151
-24 -60 25 -52
2 U1
-2 -61 12 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
45097.7 0
0
29
2 1 2 0 0 4096 0 5 4 0 0 2
655 321
655 364
2 2 2 0 0 0 0 6 5 0 0 2
655 295
655 321
1 0 3 0 0 0 0 5 0 0 4 2
635 321
635 321
13 0 3 0 0 12416 0 7 0 0 0 4
263 455
253 455
253 321
640 321
1 0 4 0 0 4096 0 11 0 0 20 2
329 193
368 193
2 0 2 0 0 4096 0 11 0 0 16 2
329 202
400 202
3 0 2 0 0 0 0 11 0 0 16 2
329 211
400 211
5 0 2 0 0 0 0 11 0 0 16 2
329 229
400 229
6 0 4 0 0 0 0 11 0 0 20 2
329 238
368 238
7 0 4 0 0 0 0 11 0 0 20 2
329 247
368 247
8 0 2 0 0 0 0 11 0 0 16 2
329 256
400 256
4 0 4 0 0 0 0 11 0 0 20 2
329 220
368 220
4 0 2 0 0 4096 0 7 0 0 16 2
327 428
400 428
6 0 2 0 0 0 0 7 0 0 16 2
327 446
400 446
7 0 2 0 0 0 0 7 0 0 16 2
327 455
400 455
1 8 2 0 0 4224 0 8 7 0 0 3
400 108
400 464
327 464
3 0 4 0 0 4096 0 7 0 0 20 2
327 419
368 419
2 0 4 0 0 0 0 7 0 0 20 2
327 410
368 410
1 0 4 0 0 0 0 7 0 0 20 2
327 401
368 401
1 5 4 0 0 4224 0 10 7 0 0 3
368 110
368 437
327 437
13 1 5 0 0 12416 0 11 6 0 0 4
265 247
253 247
253 295
635 295
0 9 2 0 0 0 0 0 7 28 0 3
234 193
234 401
257 401
0 12 6 0 0 4096 0 0 7 26 0 3
208 328
208 428
263 428
0 11 7 0 0 4224 0 0 7 27 0 3
201 313
201 419
263 419
0 10 8 0 0 4224 0 0 7 29 0 3
197 298
197 410
263 410
1 12 6 0 0 8320 0 3 11 0 0 4
183 328
208 328
208 220
265 220
1 11 7 0 0 0 0 2 11 0 0 4
183 313
203 313
203 211
265 211
1 9 2 0 0 128 0 9 11 0 0 3
234 111
234 193
259 193
1 10 8 0 0 128 0 1 11 0 0 4
183 298
198 298
198 202
265 202
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
3
13 Logic Switch~
5 397 300 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3857 0 0
2
5.90077e-315 0
0
7 Ground~
168 622 334 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7125 0 0
2
5.90077e-315 0
0
4 LED~
171 622 310 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
1 S
27 -10 34 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3641 0 0
2
5.90077e-315 0
0
2
1 1 3 0 0 8320 0 1 3 0 0 2
409 300
622 300
2 1 2 0 0 4224 0 3 2 0 0 2
622 320
622 328
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 61
913 317 1006 441
923 325 995 421
61 A  B  | S 
0  0  | X   
0  1  | 0  
1  0  | 1  
1  1  | 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 281
733 123 1250 307
743 131 1239 275
281 Entradas:
A: sensor rua A, (0: sem carros transitando, 1: carros 
transitando)
B: sensor rua B, (0: sem carros transitando, 1: carros 
transitantdo)

Sa�das:
S: controle dos sem�foros, (0: sem�foro 1 vermelho, sem�foro 2 
verde, 1: sem�foro 1 verde, sem�foro 2 vermelho)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

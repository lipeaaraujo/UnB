CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 316 303 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
45067.5 0
0
13 Logic Switch~
5 317 263 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
45067.5 1
0
13 Logic Switch~
5 316 222 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
45067.5 2
0
13 Logic Switch~
5 316 185 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
45067.5 3
0
9 3-In AND~
219 404 261 0 4 22
0 7 8 6 4
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
8157 0 0
2
45067.5 4
0
8 2-In OR~
219 465 231 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5572 0 0
2
45067.5 5
0
7 Ground~
168 529 298 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
45067.5 6
0
4 LED~
171 529 266 0 2 2
10 3 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
45067.5 7
0
7
3 1 3 0 0 4224 0 6 8 0 0 3
498 231
529 231
529 256
4 2 4 0 0 12416 0 5 6 0 0 4
425 261
429 261
429 240
452 240
1 1 5 0 0 4224 0 4 6 0 0 4
328 185
398 185
398 222
452 222
1 3 6 0 0 8320 0 1 5 0 0 4
328 303
357 303
357 270
380 270
1 1 7 0 0 8320 0 3 5 0 0 4
328 222
356 222
356 252
380 252
1 2 8 0 0 8320 0 2 5 0 0 3
329 263
329 261
380 261
2 1 2 0 0 4224 0 8 7 0 0 4
529 276
529 320
529 320
529 292
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 207
616 81 1069 245
626 89 1058 217
207 Entradas:
A, B, C e D. S�o os bits que representam, na ordem do 
mais significativo para o menos significativo, o valor 
da tens�o da bateria.

Sa�das:
S: lamp�da do painel, (0: desligada, 1: ligada)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 287
741 251 882 595
751 259 871 531
287 A  B  C  D  | S
0  0  0  0  | 0
0  0  0  1  | 0
0  0  1  0  | 0
0  0  1  1  | 0
0  1  0  0  | 0
0  1  0  1  | 0
0  1  1  0  | 0
0  1  1  1  | 1
1  0  0  0  | 1
1  0  0  1  | 1
1  0  1  0  | 1
1  0  1  1  | 1
1  1  0  0  | 1
1  1  0  1  | 1
1  1  1  0  | 1
1  1  1  1  | 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

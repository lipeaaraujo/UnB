CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
4
13 Logic Switch~
5 398 302 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 M
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5789 0 0
2
45062.9 0
0
7 Ground~
168 622 334 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7328 0 0
2
45062.9 1
0
4 LED~
171 622 310 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
5 ABRIR
14 -10 49 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4799 0 0
2
45062.9 2
0
5 4049~
219 489 301 0 2 22
0 4 3
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
9196 0 0
2
45062.9 3
0
3
2 1 2 0 0 4224 0 3 2 0 0 2
622 320
622 328
2 1 3 0 0 8320 0 4 3 0 0 3
510 301
510 300
622 300
1 1 4 0 0 8320 0 1 4 0 0 3
410 302
410 301
474 301
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 288
891 272 1040 616
901 280 1029 552
288 A  B  C  D  | S1
0  0  0  0  | X
0  0  0  1  | 1
0  0  1  0  | 1
0  0  1  1  | X
0  1  0  0  | 1
0  1  0  1  | X
0  1  1  0  | X
0  1  1  1  | X
1  0  0  0  | 0
1  0  0  1  | 0
1  0  1  0  | 0
1  0  1  1  | X
1  1  0  0  | 0
1  1  0  1  | X
1  1  1  0  | X
1  1  1  1  | X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 351
713 67 1262 251
723 75 1251 219
351 Entradas:
M: movimento do elevador (0: parado, 1: em movimento)
F1: sensor andar 1, (0: elevador presente, 1: elevador presente)
F2: sensor andar 2, (0: elevador presente, 1: elevador presente)
F3: sensor andar 3, (0: elevador presente, 1: elevador presente)

Sa�das:
ABRIR: sinal da porta, (0: sinal para porta, 1: sinal para a porta 
abrir)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

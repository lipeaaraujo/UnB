CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 290 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 173 541 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 173 503 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 173 464 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90077e-315 0
0
13 Logic Switch~
5 174 426 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90077e-315 0
0
4 LED~
171 499 375 0 2 2
10 4 2
0
0 0 880 90
4 LED1
-12 -21 16 -13
2 B1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3536 0 0
2
5.90077e-315 0
0
9 Inverter~
13 316 292 0 2 22
0 7 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
4597 0 0
2
5.90077e-315 0
0
9 Inverter~
13 316 255 0 2 22
0 8 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3835 0 0
2
5.90077e-315 0
0
9 Inverter~
13 315 356 0 2 22
0 12 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3670 0 0
2
5.90077e-315 0
0
9 Inverter~
13 314 400 0 2 22
0 11 10
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
5616 0 0
2
5.90077e-315 0
0
4 LED~
171 499 274 0 2 2
10 3 2
0
0 0 880 90
4 LED1
-12 -21 16 -13
2 B2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9323 0 0
2
5.90077e-315 0
0
7 Ground~
168 558 411 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
5.90077e-315 0
0
9 2-In AND~
219 394 376 0 3 22
0 9 10 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3108 0 0
2
5.90077e-315 0
0
9 2-In AND~
219 395 275 0 3 22
0 6 5 3
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4299 0 0
2
5.90077e-315 0
0
12
2 0 2 0 0 4096 0 5 0 0 2 2
512 376
558 376
2 1 2 0 0 8320 0 10 11 0 0 3
512 275
558 275
558 405
3 1 3 0 0 4224 0 13 10 0 0 2
416 275
492 275
3 1 4 0 0 4224 0 12 5 0 0 2
415 376
492 376
2 2 5 0 0 12416 0 6 13 0 0 4
337 292
353 292
353 284
371 284
2 1 6 0 0 12416 0 7 13 0 0 4
337 255
353 255
353 266
371 266
1 1 7 0 0 8320 0 1 6 0 0 4
185 541
251 541
251 292
301 292
1 1 8 0 0 8320 0 3 7 0 0 4
185 464
217 464
217 255
301 255
2 1 9 0 0 4224 0 8 12 0 0 4
336 356
353 356
353 367
370 367
2 2 10 0 0 4224 0 9 12 0 0 4
335 400
353 400
353 385
370 385
1 1 11 0 0 8320 0 2 9 0 0 4
185 503
234 503
234 400
299 400
1 1 12 0 0 12416 0 4 8 0 0 4
186 426
201 426
201 356
300 356
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 339
722 395 895 739
732 403 884 675
339 S1 S2 S3 S4 | B1 B2
0  0  0  0  | 1  1
0  0  0  1  | 1  0
0  0  1  0  | 0  1
0  0  1  1  | 0  0
0  1  0  0  | 1  0
0  1  0  1  | 1  0
0  1  1  0  | 0  0
0  1  1  1  | 0  0
1  0  0  0  | 0  1
1  0  0  1  | 0  0
1  0  1  0  | 0  1
1  0  1  1  | 0  0
1  1  0  0  | 0  0
1  1  0  1  | 0  0
1  1  1  0  | 0  0
1  1  1  1  | 0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 472
647 136 1116 440
657 144 1105 384
472 Entradas:
S1: sensor de n�vel baixo do T1
(0: n�vel n�o baixo, 1: n�vel baixo)
S2: sensor de n�vel baixo do T2
(0: n�vel n�o baixo, 1: n�vel baixo)
S3: sensor de n�vel m�ximo do T2
(0: n�vel m�ximo n�o atingido, 1: n�vel m�ximo atingido)
S4: sensor de n�vel m�ximo do T3
(0: n�vel m�ximo n�o atingido, 1: n�vel m�ximo atingido)

Sa�das:
B1: bomba do tanque T1
(0: bomba desligada, 1: bomba ligada)
B2: bomba do tanque T2
(0: bomba desligada, 1: bomba ligada)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 192
319 443 716 527
329 451 705 515
192 A bomba B1 ficar� ligada quando o tanque T1 n�o
estiver vazio e o tanque T2 n�o estiver cheio.
A bomba B2 ficar� ligada quando o tanque T2 n�o
estiver vazio e o tanque T3 n�o estiver cheio.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 339 369 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90083e-315 0
0
13 Logic Switch~
5 143 284 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90083e-315 0
0
13 Logic Switch~
5 298 158 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.90083e-315 0
0
13 Logic Switch~
5 318 158 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.90083e-315 0
0
4 LED~
171 621 357 0 2 2
10 8 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8157 0 0
2
5.90083e-315 0
0
4 LED~
171 622 469 0 2 2
10 5 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5572 0 0
2
5.90083e-315 0
0
4 LED~
171 622 430 0 2 2
10 6 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8901 0 0
2
5.90083e-315 0
0
4 LED~
171 622 394 0 2 2
10 7 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
5.90083e-315 0
0
7 Ground~
168 435 170 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.90083e-315 0
0
2 +V
167 457 173 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.90083e-315 0
0
7 74LS194
49 389 333 0 14 29
0 11 10 9 2 4 3 4 2 4
2 8 7 6 5
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3472 0 0
2
5.90083e-315 0
0
18
1 6 3 0 0 0 0 1 11 0 0 2
351 369
351 369
5 0 4 0 0 12288 0 11 0 0 17 4
357 351
347 351
347 268
457 268
2 0 2 0 0 12416 0 6 0 0 15 4
622 479
701 479
701 224
435 224
2 0 2 0 0 0 0 7 0 0 15 4
622 440
691 440
691 234
435 234
2 0 2 0 0 0 0 8 0 0 15 4
622 404
681 404
681 244
435 244
2 0 2 0 0 0 0 5 0 0 15 4
621 367
671 367
671 253
435 253
4 0 2 0 0 0 0 11 0 0 15 3
357 342
357 263
435 263
14 1 5 0 0 4224 0 11 6 0 0 4
421 369
587 369
587 459
622 459
13 1 6 0 0 4224 0 11 7 0 0 4
421 360
595 360
595 420
622 420
12 1 7 0 0 4224 0 11 8 0 0 4
421 351
603 351
603 384
622 384
11 1 8 0 0 4224 0 11 5 0 0 3
421 342
621 342
621 347
1 3 9 0 0 4224 0 4 11 0 0 3
318 170
318 324
357 324
1 2 10 0 0 4224 0 3 11 0 0 3
298 170
298 315
357 315
0 10 2 0 0 0 0 0 11 15 0 3
435 306
435 324
421 324
1 8 2 0 0 0 0 9 11 0 0 3
435 178
435 306
421 306
9 0 4 0 0 0 0 11 0 0 17 3
421 315
457 315
457 296
1 7 4 0 0 4224 0 10 11 0 0 3
457 182
457 297
421 297
1 1 11 0 0 4224 0 11 2 0 0 3
357 297
143 297
143 296
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 0 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
86 C:\Users\felip\OneDrive\�rea de Trabalho\UNB\3� Semestre\TED\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 48 181 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21488 0
2 5V
-6 -16 8 -8
2 S7
-30 -5 -16 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
631 0 0
2
45097.7 4
0
13 Logic Switch~
5 50 155 0 1 11
0 8
0
0 0 21488 0
2 0V
-6 -16 8 -8
2 S6
-30 -5 -16 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9466 0 0
2
45097.7 3
0
13 Logic Switch~
5 49 130 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21488 0
2 5V
-6 -16 8 -8
2 S5
-30 -4 -16 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3266 0 0
2
45097.7 2
0
13 Logic Switch~
5 48 105 0 1 11
0 4
0
0 0 21488 0
2 0V
-6 -16 8 -8
2 S4
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7693 0 0
2
45097.7 1
0
9 Inverter~
13 168 72 0 2 22
0 4 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3723 0 0
2
45097.8 0
0
4 LED~
171 675 216 0 1 2
10 10
0
0 0 352 90
2 S0
-20 4 -6 12
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3440 0 0
2
45097.7 0
0
4 LED~
171 675 194 0 1 2
10 13
0
0 0 352 90
2 S1
-20 5 -6 13
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6263 0 0
2
45097.7 0
0
4 LED~
171 676 173 0 1 2
10 6
0
0 0 352 90
2 S2
-21 5 -7 13
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4900 0 0
2
45097.7 0
0
4 LED~
171 676 152 0 1 2
10 18
0
0 0 352 90
2 S3
-20 5 -6 13
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8783 0 0
2
45097.7 0
0
7 74LS151
20 237 746 0 14 29
0 3 3 3 3 3 3 3 3 5
9 8 7 12 21
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
3221 0 0
2
45097.7 2
0
7 74LS151
20 237 861 0 14 29
0 2 2 2 2 2 2 2 2 4
9 8 7 11 22
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
3215 0 0
2
45097.7 1
0
8 2-In OR~
219 424 799 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7903 0 0
2
45097.7 0
0
7 74LS151
20 238 530 0 14 29
0 2 2 2 2 3 3 3 3 5
9 8 7 15 23
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
7121 0 0
2
45097.7 2
0
7 74LS151
20 238 645 0 14 29
0 3 3 3 3 2 2 2 2 4
9 8 7 14 24
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
4484 0 0
2
45097.7 1
0
8 2-In OR~
219 425 583 0 3 22
0 15 14 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5996 0 0
2
45097.7 0
0
7 74LS151
20 239 315 0 14 29
0 2 2 3 3 3 3 2 2 5
9 8 7 17 25
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
7804 0 0
2
45097.7 2
0
7 74LS151
20 239 430 0 14 29
0 2 2 3 3 3 3 2 2 4
9 8 7 16 26
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
5523 0 0
2
45097.7 1
0
8 2-In OR~
219 426 368 0 3 22
0 17 16 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3330 0 0
2
45097.7 0
0
8 2-In OR~
219 426 153 0 3 22
0 20 19 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3465 0 0
2
45097.7 0
0
7 74LS151
20 239 215 0 14 29
0 2 3 3 2 2 3 3 2 4
9 8 7 19 27
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
8396 0 0
2
45097.7 6
0
7 74LS151
20 239 100 0 14 29
0 2 3 3 2 2 3 3 2 5
9 8 7 20 28
0
0 0 4336 512
7 74LS151
-24 -60 25 -52
0
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
3685 0 0
2
45097.7 5
0
2 +V
167 331 26 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7849 0 0
2
45097.7 0
0
7 Ground~
168 357 31 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6343 0 0
2
45097.7 0
0
113
2 0 0 0 0 0 0 9 0 0 71 3
689 153
689 52
357 52
2 2 0 0 0 0 0 8 9 0 0 2
689 174
689 153
2 2 0 0 0 0 0 7 8 0 0 3
688 195
689 195
689 174
2 2 0 0 0 0 0 6 7 0 0 2
688 217
688 195
1 0 2 0 0 4096 0 21 0 0 71 2
277 73
357 73
2 0 3 0 0 4096 0 21 0 0 65 2
277 82
331 82
3 0 3 0 0 0 0 21 0 0 65 2
277 91
331 91
4 0 2 0 0 0 0 21 0 0 71 2
277 100
357 100
5 0 2 0 0 0 0 21 0 0 71 2
277 109
357 109
6 0 3 0 0 0 0 21 0 0 65 2
277 118
331 118
7 0 3 0 0 0 0 21 0 0 65 2
277 127
331 127
8 0 2 0 0 0 0 21 0 0 71 2
277 136
357 136
1 0 2 0 0 0 0 20 0 0 71 2
277 188
357 188
2 0 3 0 0 0 0 20 0 0 65 2
277 197
331 197
3 0 3 0 0 0 0 20 0 0 65 2
277 206
331 206
4 0 2 0 0 0 0 20 0 0 71 2
277 215
357 215
5 0 2 0 0 0 0 20 0 0 71 2
277 224
357 224
6 0 3 0 0 0 0 20 0 0 65 2
277 233
331 233
7 0 3 0 0 0 0 20 0 0 65 2
277 242
331 242
8 0 2 0 0 0 0 20 0 0 71 2
277 251
357 251
0 1 4 0 0 4096 0 0 5 23 0 3
146 105
146 72
153 72
9 2 5 0 0 8192 0 21 5 0 0 3
207 73
207 72
189 72
1 0 4 0 0 4096 0 4 0 0 96 3
60 105
146 105
146 188
1 0 2 0 0 4096 0 11 0 0 71 2
275 834
357 834
2 0 2 0 0 0 0 11 0 0 71 2
275 843
357 843
1 0 2 0 0 0 0 16 0 0 71 2
277 288
357 288
2 0 2 0 0 0 0 16 0 0 71 2
277 297
357 297
3 0 3 0 0 0 0 16 0 0 65 2
277 306
331 306
4 0 3 0 0 0 0 16 0 0 65 2
277 315
331 315
5 0 3 0 0 0 0 16 0 0 65 2
277 324
331 324
6 0 3 0 0 0 0 16 0 0 65 2
277 333
331 333
7 0 2 0 0 0 0 16 0 0 71 2
277 342
357 342
8 0 2 0 0 0 0 16 0 0 71 2
277 351
357 351
1 0 2 0 0 0 0 17 0 0 71 2
277 403
357 403
2 0 2 0 0 0 0 17 0 0 71 2
277 412
357 412
3 0 3 0 0 0 0 17 0 0 65 2
277 421
331 421
4 0 3 0 0 0 0 17 0 0 65 2
277 430
331 430
5 0 3 0 0 0 0 17 0 0 65 2
277 439
331 439
6 0 3 0 0 0 0 17 0 0 65 2
277 448
331 448
7 0 2 0 0 0 0 17 0 0 71 2
277 457
357 457
8 0 2 0 0 0 0 17 0 0 71 2
277 466
357 466
1 0 2 0 0 0 0 13 0 0 71 2
276 503
357 503
2 0 2 0 0 0 0 13 0 0 71 2
276 512
357 512
3 0 2 0 0 0 0 13 0 0 71 2
276 521
357 521
4 0 2 0 0 0 0 13 0 0 71 2
276 530
357 530
5 0 3 0 0 4096 0 13 0 0 65 2
276 539
331 539
6 0 3 0 0 0 0 13 0 0 65 2
276 548
331 548
7 0 3 0 0 0 0 13 0 0 65 2
276 557
331 557
8 0 3 0 0 0 0 13 0 0 65 2
276 566
331 566
1 0 3 0 0 0 0 14 0 0 65 2
276 618
331 618
2 0 3 0 0 0 0 14 0 0 65 2
276 627
331 627
3 0 3 0 0 0 0 14 0 0 65 2
276 636
331 636
4 0 3 0 0 0 0 14 0 0 65 2
276 645
331 645
5 0 2 0 0 0 0 14 0 0 71 2
276 654
357 654
6 0 2 0 0 0 0 14 0 0 71 2
276 663
357 663
7 0 2 0 0 0 0 14 0 0 71 2
276 672
357 672
8 0 2 0 0 0 0 14 0 0 71 2
276 681
357 681
1 0 3 0 0 4096 0 10 0 0 65 2
275 719
331 719
2 0 3 0 0 0 0 10 0 0 65 2
275 728
331 728
3 0 3 0 0 0 0 10 0 0 65 2
275 737
331 737
4 0 3 0 0 0 0 10 0 0 65 2
275 746
331 746
5 0 3 0 0 0 0 10 0 0 65 2
275 755
331 755
6 0 3 0 0 0 0 10 0 0 65 2
275 764
331 764
7 0 3 0 0 0 0 10 0 0 65 2
275 773
331 773
1 8 3 0 0 4224 0 22 10 0 0 3
331 35
331 782
275 782
3 0 2 0 0 0 0 11 0 0 71 2
275 852
357 852
4 0 2 0 0 0 0 11 0 0 71 2
275 861
357 861
5 0 2 0 0 0 0 11 0 0 71 2
275 870
357 870
6 0 2 0 0 0 0 11 0 0 71 2
275 879
357 879
7 0 2 0 0 0 0 11 0 0 71 2
275 888
357 888
1 8 2 0 0 4224 0 23 11 0 0 3
357 39
357 897
275 897
3 1 6 0 0 8320 0 18 8 0 0 4
459 368
577 368
577 174
669 174
12 0 7 0 0 4096 0 16 0 0 78 2
213 315
155 315
12 0 7 0 0 0 0 17 0 0 78 2
213 430
155 430
12 0 7 0 0 0 0 13 0 0 78 2
212 530
155 530
12 0 7 0 0 0 0 14 0 0 78 2
212 645
155 645
12 0 7 0 0 0 0 10 0 0 78 2
211 746
155 746
0 12 7 0 0 4224 0 0 11 111 0 3
155 212
155 861
211 861
11 0 8 0 0 4096 0 16 0 0 84 2
213 306
163 306
11 0 8 0 0 0 0 17 0 0 84 2
213 421
163 421
11 0 8 0 0 0 0 13 0 0 84 2
212 521
163 521
11 0 8 0 0 0 0 14 0 0 84 2
212 636
163 636
11 0 8 0 0 0 0 10 0 0 84 2
211 737
163 737
0 11 8 0 0 4224 0 0 11 112 0 3
163 205
163 852
211 852
10 0 9 0 0 4096 0 14 0 0 90 2
212 627
170 627
10 0 9 0 0 4096 0 16 0 0 90 2
213 297
170 297
10 0 9 0 0 0 0 17 0 0 90 2
213 412
170 412
10 0 9 0 0 0 0 13 0 0 90 2
212 512
170 512
10 0 9 0 0 0 0 10 0 0 90 2
211 728
170 728
0 10 9 0 0 4224 0 0 11 113 0 3
170 195
170 843
211 843
9 9 5 0 0 8320 0 13 10 0 0 3
206 503
205 503
205 719
9 9 5 0 0 0 0 16 13 0 0 3
207 288
206 288
206 503
9 9 5 0 0 0 0 21 16 0 0 2
207 73
207 288
9 0 4 0 0 0 0 17 0 0 96 2
207 403
146 403
9 0 4 0 0 0 0 14 0 0 96 2
206 618
146 618
9 9 4 0 0 8320 0 20 11 0 0 4
207 188
146 188
146 834
205 834
3 1 10 0 0 8320 0 12 6 0 0 4
457 799
627 799
627 217
668 217
13 2 11 0 0 8320 0 11 12 0 0 5
211 888
211 800
403 800
403 808
411 808
13 1 12 0 0 8320 0 10 12 0 0 5
211 773
211 795
403 795
403 790
411 790
3 1 13 0 0 8320 0 15 7 0 0 4
458 583
602 583
602 195
668 195
13 2 14 0 0 8320 0 14 15 0 0 5
212 672
212 584
404 584
404 592
412 592
13 1 15 0 0 8320 0 13 15 0 0 5
212 557
212 579
404 579
404 574
412 574
13 2 16 0 0 8320 0 17 18 0 0 5
213 457
213 369
405 369
405 377
413 377
13 1 17 0 0 8320 0 16 18 0 0 5
213 342
213 364
405 364
405 359
413 359
3 1 18 0 0 4224 0 19 9 0 0 2
459 153
669 153
13 2 19 0 0 8320 0 20 19 0 0 5
213 242
213 154
405 154
405 162
413 162
13 1 20 0 0 8320 0 21 19 0 0 5
213 127
213 149
405 149
405 144
413 144
0 12 7 0 0 0 0 0 21 111 0 3
154 181
154 100
213 100
0 11 8 0 0 0 0 0 21 112 0 3
163 155
163 91
213 91
0 10 9 0 0 0 0 0 21 113 0 3
170 130
170 82
213 82
1 12 7 0 0 0 0 1 20 0 0 4
60 181
155 181
155 215
213 215
1 11 8 0 0 0 0 2 20 0 0 4
62 155
163 155
163 206
213 206
1 10 9 0 0 0 0 3 20 0 0 4
61 130
170 130
170 197
213 197
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
